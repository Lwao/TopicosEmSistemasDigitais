library verilog;
use verilog.vl_types.all;
entity onehot_fsm_vlg_vec_tst is
end onehot_fsm_vlg_vec_tst;
