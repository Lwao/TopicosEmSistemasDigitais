library verilog;
use verilog.vl_types.all;
entity seven_segment_decoder_vlg_sample_tst is
    port(
        SW              : in     vl_logic_vector(17 downto 0);
        sampler_tx      : out    vl_logic
    );
end seven_segment_decoder_vlg_sample_tst;
