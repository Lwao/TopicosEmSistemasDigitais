library verilog;
use verilog.vl_types.all;
entity Memento_vlg_vec_tst is
end Memento_vlg_vec_tst;
