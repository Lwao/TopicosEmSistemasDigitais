library verilog;
use verilog.vl_types.all;
entity buffered_mux_vlg_vec_tst is
end buffered_mux_vlg_vec_tst;
