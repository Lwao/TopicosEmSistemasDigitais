library verilog;
use verilog.vl_types.all;
entity counter3_vlg_vec_tst is
end counter3_vlg_vec_tst;
