LIBRARY ieee;
USE ieee.std_logic_1164.all;

PACKAGE MementoComponents IS

	COMPONENT AddSub is
		GENERIC (n : INTEGER := 16);
		PORT(
			 X, Y: IN STD_LOGIC_VECTOR (n-1 DOWNTO 0);
			 MUX: IN STD_LOGIC;
			 Z: OUT STD_LOGIC_VECTOR (n-1 DOWNTO 0);
			 C, V: OUT STD_LOGIC
			);
	END COMPONENT AddSub;
	
	COMPONENT UpCounter IS
		PORT (
			Clear, Clock : IN STD_LOGIC;
			Q : OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
		);
	END COMPONENT UpCounter;
	
	COMPONENT Decoder3to8 IS
		PORT (
			W : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
			En : IN STD_LOGIC;
			Y : OUT STD_LOGIC_VECTOR(0 TO 7)
		);
	END COMPONENT Decoder3to8;
	
	COMPONENT MultiplexerN IS
		GENERIC (n : INTEGER := 16);
		PORT (
			R0, R1, R2, R3, R4, R5, R6, R7, DIN, G: IN STD_LOGIC_VECTOR(n-1 DOWNTO 0);
			sel: IN STD_LOGIC_VECTOR(9 DOWNTO 0);
			ena: IN STD_LOGIC;
			y: OUT STD_LOGIC_VECTOR(n-1 DOWNTO 0)
		);
	END COMPONENT MultiplexerN;
	
	COMPONENT RegisterN IS
		GENERIC (n : INTEGER := 16);
		PORT (
			R : IN STD_LOGIC_VECTOR(n-1 DOWNTO 0);
			Rin, Clock : IN STD_LOGIC;
			Q : BUFFER STD_LOGIC_VECTOR(n-1 DOWNTO 0)
		);
	END COMPONENT RegisterN;


END PACKAGE MementoComponents;