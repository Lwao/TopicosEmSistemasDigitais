library verilog;
use verilog.vl_types.all;
entity dff1_vlg_vec_tst is
end dff1_vlg_vec_tst;
